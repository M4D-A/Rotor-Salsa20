module double_round_tb;

// Clock and step counter
parameter CLKp = 10;
reg clk = 1'b0;
reg [31:0] ctr = 32'b0;

always begin
	#(CLKp/2) clk = !clk;
end

// unit test data and control
reg [511:0] unit_data [0:15];
reg [31:0] correct_ctr = 32'b0;
reg test_passed = 1'b0;
wire correct;

// Testbench block IO
reg [511:0] in;
wire [511:0] out;

// Success Condition
assign correct = (out == unit_data[ctr]) ? 1'b1 : 1'b0;

// Initialize unit test data
initial begin
    unit_data[00][511:256] <= 256'hAE2F43E8_2BEB539C_A50ED7EF_F7D2876_B0000000_00CD7B55_408D4BC9_0E48046A5;
    unit_data[00][255:000] <= 256'h77EF56DF_6FBBF7AB_07E6DBF6_3F0E2B1_A8025E49_5AD442EB_C7767D27_3ABAA7A0C;
    unit_data[01][511:256] <= 256'h4A49D6B2_A437B0E5_52C6BD8F_937772C_5C0D9B0A_C09995F9_90A95F47_F21AB7807;
    unit_data[01][255:000] <= 256'h0A88D59F_19059A54_E5ED16F0_4C70F4B_AC74DFBC_B5F6ED64_FF8DBB00_0567ADEF9;
    unit_data[02][511:256] <= 256'h5FF3F20B_E41B15F5_65C72C3C_36414E4_6687E956_DCDA539E_62652B95_C41E3AFB4;
    unit_data[02][255:000] <= 256'h8086DF19_905DA17D_70911C4F_254AE9D_26CF75DF_041AB31A_10846A22_7C5E3985D;
    unit_data[03][511:256] <= 256'h4363666C_B93AFD62_EB3EF7AB_DE83EAB_78C3E508_D784626C_AEBFB348_32ADEE328;
    unit_data[03][255:000] <= 256'h165AEC92_9817998B_319DDAA8_67FA0DE_2BE4420D_F3D78F00_4CCE66F8_2D730A6EA;
    unit_data[04][511:256] <= 256'h0D682289_6A7E3311_E6E44229_40FBAAF_E083CD06_D6B1AF19_B83A3348_1A3AC837B;
    unit_data[04][255:000] <= 256'h9E65C005_9572F116_8972CBC1_AB91BB4_3E506DBF_F26BF138_B177D494_17E07FB13;
    unit_data[05][511:256] <= 256'h63B5709F_B3D2B717_3E22CF63_A6122B8_B61E2466_C4052D12_B716B781_00C2A0FAA;
    unit_data[05][255:000] <= 256'h28DEC5CE_3512060F_1BEBE8B2_3339182_2830E835_52BE4976_2F1210C2_798D55F0B;
    unit_data[06][511:256] <= 256'h99840033_9A419D77_B9CF2478_0105BB4_D54E30D6_274630E3_643CB2B2_1A8DA996F;
    unit_data[06][255:000] <= 256'h066E25DE_ADB3BAAD_D8B77914_7CED25B_9FED35B0_3D66C323_D17397DF_5E3B895EB;
    unit_data[07][511:256] <= 256'h4914F6DE_AD3287CD_B0029493_A9574C2_80149471_A92695A7_002DEFE1_A8D1C8458;
    unit_data[07][255:000] <= 256'h0720C75D_B552E970_248F3815_55DC0E4_519CB95A_750E29A1_BD1BC0AD_5FA061BCB;
    unit_data[08][511:256] <= 256'hB7F159DF_21398D45_C7542512_0E066C4_543FEC8F_297C8488_BA29089D_ED1FD6686;
    unit_data[08][255:000] <= 256'h539F975C_78B37A7B_9367769F_99550E1_E86E7DB7_47E053A3_319B0476_2A1274998;
    unit_data[09][511:256] <= 256'h7A974624_51297A9C_F6A6C21B_AFE3AD7_0EB9D213_A10CE816_0D0A04F6_047AAAE44;
    unit_data[09][255:000] <= 256'h9F9C3B2F_01C95005_CD15C6AF_BEE974E_5ED3640D_EDE4CDC4_CBC6FC1B_BBBAB9E7C;
    unit_data[10][511:256] <= 256'h8ABC872B_42814A1B_DE58865F_321A3BA_5DC5C6F8_7408757D_B0D16D13_57C2C8C0E;
    unit_data[10][255:000] <= 256'h76B0AFAB_45BEC005_FA0ACDFB_94BA955_D246092F_B56068CB_B92B00E7_0C37DB471;
    unit_data[11][511:256] <= 256'hCAC64FE0_413304D6_35FE373B_BE72CE9_227319F5_51E7CFB9_4640CED8_62478044B;
    unit_data[11][255:000] <= 256'h554737FA_37FF3150_FC6DE923_926BCF8_FAA6BB36_01A6F4FB_AAAD0C3C_97B887065;
    unit_data[12][511:256] <= 256'h3F2617C7_C5ACAB0F_F72CCB6A_F86908E_4866D242_04503587_B461FBBB_07CC0C609;
    unit_data[12][255:000] <= 256'h5172A009_DFAC9EDE_CED4A2BE_8828523_0AEE197D_FDAC5A9B_E177A522_F8E31F32E;
    unit_data[13][511:256] <= 256'hECDA2537_511F3BE7_20BC4454_C319D5E_D9A622A3_F3731174_8A5A60E8_A83EBFBDF;
    unit_data[13][255:000] <= 256'h9CD15ECE_B4A9293F_50334019_9457F15_C39FE7DA_339F925B_692F9CE5_ACD57FFDA;
    unit_data[14][511:256] <= 256'h6F0012D4_A6F57D75_CE873347_5CB1A30_92208A5C_67350D0C_17A05B79_5E569A35E;
    unit_data[14][255:000] <= 256'hE19B9C05_26E3CEA0_F4A9F4C3_41E9B39_BEBE3871_AB86A630_85767FEC_AFC42D918;
    unit_data[15][511:256] <= 256'hC2327B61_1DE9EE83_17DCEEFB_02001B9_E2AC091B_07892A99_A7D10A8C_4A4F7EDB6;
    unit_data[15][255:000] <= 256'h30DE3E65_63D175C1_4B19F2F0_CD5371A_22C68D95_67FC4655_E185DB95_AF9D82094;
end

// Initialize testbenched block inputs
initial begin 
    in[255:000] <= 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_deadbeef;
    in[512:256] <= 256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_feedface;
end

// Testbench block control
always @(posedge clk) begin
    in <= out; // Forward output to input

    correct_ctr <= (correct == 1'b1) ? correct_ctr + 1'b1 : correct_ctr;
    test_passed <= (correct_ctr == 31'd16) ? 1'b1 : 1'b0;
    if(ctr == 31'd16) begin
        if(correct_ctr == 16) begin
            $display("TEST PASSED: ", correct_ctr," /16 correct results");
        end 
        else begin
            $display("TEST FAILED", correct_ctr);
        end
        $finish;
    end 

    ctr <= ctr + 1'b1;
end

double_round tb_block(
    .d_in(in),
    .d_out(out)
);

endmodule


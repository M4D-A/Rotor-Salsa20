module salsa_hash_tb;

// Clock and step counter
parameter CLKp = 10;
reg clk = 1'b0;
reg [31:0] ctr = 32'b0;

always begin
	#(CLKp/2) clk = !clk;
end

// unit test data and control
reg [511:0] unit_data [0:15];
reg [31:0] correct_ctr = 32'b0;
reg test_passed = 1'b0;
wire correct;

// Testbench block IO
reg  [255 : 0] key_in = 256'h80;
reg  [63 : 0] nonce_in = 64'h0;
reg  [63 : 0] counter_in = 64'h0;
wire [511 : 0] digest_out;

// Success Condition
assign correct = (digest_out == unit_data[ctr]) ? 1'b1 : 1'b0;

// Initialize unit test data
initial begin
    unit_data[00][511:256] <= 256'h_17A1F17E_4DAF7618_469C2AE7_832A6544_079A8DFC_E43FBDCB_C723279E_55972CB2;
    unit_data[00][255:000] <= 256'h_44689FAD_5F7A3BD2_385C7A09_E1513900_E7A6295B_47F98EEA_E3A2EC8B_DD8FBEE3;
    unit_data[01][511:256] <= 256'h_AE48E353_B2B4CD93_F7505126_F146120F_BB6E6D36_56F46926_2AD117A1_A90314CC;
    unit_data[01][255:000] <= 256'h_01208056_C3C5206B_6B81E269_466E71E9_38E5CAAB_6601E2E7_83621BEF_4EB7A28D;
    unit_data[02][511:256] <= 256'h_69D1D7F2_168DBEE3_98B461E8_74DD9F12_68530B32_50488276_7D760495_E2B14201;
    unit_data[02][255:000] <= 256'h_07844B0E_8B2B225E_8DB3D5E7_B17CE0B7_36AA701D_62000E7E_2A805E02_BC893D20;
    unit_data[03][511:256] <= 256'h_17AA1F29_73DC9FED_6A1A2EFB_F412E798_CAE11735_B68BBF8A_8EF2A76D_12CD84ED;
    unit_data[03][255:000] <= 256'h_A916624C_A7081371_3CA9903A_ED50F2AC_103EA729_54F14F7C_AED9177B_F481BE57;
    unit_data[04][511:256] <= 256'h_18B60110_D71018FB_8F0BD1D8_C72E163E_A656344B_1AB7149F_0CA4EFAC_7CF50A7C;
    unit_data[04][255:000] <= 256'h_7EAA40CE_7D65ECAE_39C0F194_E194A291_3A511FB8_ED35C638_58BD2EBA_C4118295;
    unit_data[05][511:256] <= 256'h_ED431CA4_435B2CE1_D7844058_5694305E_E7563641_B01C47C3_CEFAC600_A7319634;
    unit_data[05][255:000] <= 256'h_88E92051_B6914EEC_C7988A6D_922E7F0C_AEA80F89_2D7B1FC1_0554B853_DA739F2F;
    unit_data[06][511:256] <= 256'h_22C6BFC7_FDB7EFF4_DD828F29_AD7DDF23_7E05C79E_6A0C9293_C2FD44CE_05653E90;
    unit_data[06][255:000] <= 256'h_31B3BD32_9FF67D7F_4B64AE2C_E62F29CD_777BFE20_5A666A5F_A60D889B_BD8A049A;
    unit_data[07][511:256] <= 256'h_7784BC64_CC766AE5_364A7893_5BB132CC_55E8F108_9D080D7C_6B26A4A3_05A1EF77;
    unit_data[07][255:000] <= 256'h_536FBDA0_3399927E_13FF3596_4E35C3CD_9AD749A6_117FE7C7_83CCDD0C_FDFC6A69;
    unit_data[08][511:256] <= 256'h_E5BA89C2_C3FF926E_7EBA5235_9B8770C5_86DD1CA8_64D71B3A_3BA67355_0FAB71AC;
    unit_data[08][255:000] <= 256'h_ECF3AF59_2951CD70_82DFE111_16244F76_5EDB2789_427F2B25_CBDBA4A3_42DEA25C;
    unit_data[09][511:256] <= 256'h_BF03E4EA_8029D4D7_520C1485_117D2EDF_ECAF9A9A_31E806B5_9FBF79FB_A1F38B2B;
    unit_data[09][255:000] <= 256'h_14CD79CA_44D17454_7C51EBFC_F4EADF3E_D71EF630_FAC686A3_93AFFA0B_34CF3A56;
    unit_data[10][511:256] <= 256'h_3F66CB9F_B9B46A77_BEF306F6_09C1FB26_8E4F88E0_8DA91BC2_109DD9FD_7EC50227;
    unit_data[10][255:000] <= 256'h_009A0D71_FDAA29FC_58E8C029_9BED3E91_96FCCBBC_FD04F4CF_0D52C4D1_132CFC26;
    unit_data[11][511:256] <= 256'h_F356CFAF_ABDB18DB_8D95EBA5_E029DE4F_728C4BCB_0B6EEBD3_F2AB4459_AE36548F;
    unit_data[11][255:000] <= 256'h_6051D348_A9197DC9_6135CCBC_EA7910BA_E8050BB8_80B5F4AE_121E51D6_C73EB7EF;
    unit_data[12][511:256] <= 256'h_154EDAEC_B6BE66D7_AFD1062A_705A170F_A69D24DD_CE150B3D_5C8E9E3B_5A2D3CEC;
    unit_data[12][255:000] <= 256'h_1170A6C1_392D9AB2_8C215A74_6691B999_6B8B9494_FCB51120_0CD249A9_4C3DA608;
    unit_data[13][511:256] <= 256'h_2FF8DA97_7FFEF71E_424DF028_70633B20_5266BBB8_375117A7_8E3837C2_2156BB5A;
    unit_data[13][255:000] <= 256'h_ADEC6A74_AA4BC31A_B77CF636_6B4B58E5_27DCBEA4_37EA0F58_4ED0CEEF_E51D985A;
    unit_data[14][511:256] <= 256'h_370D4BC5_921BB441_E13477F6_11E53C83_B459E1FF_A292D045_DA53E7D2_D60452A7;
    unit_data[14][255:000] <= 256'h_D0A5792E_6970D0AC_BABB7A30_F2D64C20_D1BBAD3C_28DD934E_9A236BE4_F7419864;
    unit_data[15][511:256] <= 256'h_9D34AF3A_526DDBF2_130C44EB_DA67E2B2_FACB9CAB_3FC29D81_E79630B1_F406B058;
    unit_data[15][255:000] <= 256'h_8F5559DD_10ED4848_31328466_A0972A35_9CF5A8A6_1876C198_ADCE2A4F_2FF000A0;
end

always @(posedge clk) begin
    counter_in <= counter_in + 1'b1;

    correct_ctr <= (correct == 1'b1) ? correct_ctr + 1'b1 : correct_ctr;
    test_passed <= (correct_ctr == 31'd16) ? 1'b1 : 1'b0;
    if(ctr == 31'd16) begin
        if(correct_ctr == 16) begin
            $display("TEST PASSED: ", correct_ctr," /16 correct results");
        end 
        else begin
            $display("TEST FAILED", correct_ctr);
        end
        $finish;
    end 

    ctr <= ctr + 1'b1;
end

// Instantiate the module
salsa_hash tb_block(
    .key_in(key_in),
    .nonce_in(nonce_in),
    .counter_in(counter_in),
    .digest_out(digest_out)
);

endmodule































































